`include "./ysyx22041405_alu.v"
module ysyx22041405_EXU#(parameter WIDTH = 32)(
    input [WIDTH - 1: 0] rf_rs1,
    input [WIDTH - 1: 0] rf_rs2,
    input [WIDTH - 1: 0] Imm,
    // ALU port
    output[WIDTH - 1: 0] alu_result
);
    //======================== ALU module ================================

    
endmodule //ysyx22041405_EXU
